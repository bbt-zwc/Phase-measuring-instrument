`timescale 1ns / 1ps

module tb1();

// 输入输出信号声明
reg clk_1hz;       // 1Hz输入时钟（由测试平台生成）
reg rst_n;         // 复位信号（低有效）
reg [15:0] fre;    // 频率输入（测试中动态设置）
wire led;          // LED输出（观测目标）

// 实例化被测试模块
alarm uut (
    .clk_1hz(clk_1hz),
    .rst_n(rst_n),
    .fre(fre),
    .led(led)
);

// --------------------------
// 生成1Hz时钟（周期1秒，半周期500ms）
// --------------------------
initial begin
    clk_1hz = 0;
    forever #500_000_000 clk_1hz = ~clk_1hz;  // 每500ms翻转一次（1Hz周期）
end

// --------------------------
// 复位控制与测试流程
// --------------------------
initial begin
    // 阶段1：复位有效（rst_n=0），持续2秒
    rst_n = 0;
    fre = 16'd0;  // 随意值（复位时不关心）
    #2000_000_000;  // 2秒（足够观察复位状态）
    
    // 阶段2：复位释放（rst_n=1），设置fre≤20000（16'd10000），持续3秒
    rst_n = 1;
    fre = 16'd10000;  // 10000 ≤ 20000，LED应保持0
    #3000_000_000;  // 3秒
    
    // 阶段3：设置fre>20000（16'd30000），持续3秒
    fre = 16'd30000;  // 30000 > 20000，LED应以1Hz闪烁
    #3000_000_000;  // 3秒
    
    // 测试结束
    $finish;
end


endmodule